package apb_master_pkg;

`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "defines.sv"
`include "apb_master_seq_item.sv"
`include "apb_master_sequence.sv"
`include "apb_master_sequencer.sv"
`include "apb_master_driver.sv"
`include "apb_master_active_monitor.sv"
`include "apb_master_passive_monitor.sv"
`include "apb_master_active_agent.sv"
`include "apb_master_passive_agent.sv"
`include "apb_master_subscriber.sv"
`include "apb_master_scoreboard.sv"
`include "apb_master_env.sv"
`include "apb_master_test.sv"

endpackage
